module b;
endmodule