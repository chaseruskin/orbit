architecture arch1 of ent1 is

begin
  ok <= '1';
end architecture;