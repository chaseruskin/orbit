architecture arch2 of ent1 is

begin
  ok <= '0';
end architecture;