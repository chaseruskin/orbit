module d;
endmodule