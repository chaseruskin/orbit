entity ent1 is
  port (
    ok : out bit
  );
end entity;