module a;
endmodule