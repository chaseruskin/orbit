module top(a, b, c); 
    assign a = 1;
endmodule