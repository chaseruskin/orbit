module c;
endmodule