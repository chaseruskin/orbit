module top
    (a, b, c); 

    import ComplexPkg::*;
    
    assign a = 1;


endmodule