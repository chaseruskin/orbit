module hard timeunit 10ns / 1ns; (input clk);

endmodule: hard