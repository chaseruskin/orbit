module packer #(
    int[3:0][3:0] grid[10][1:9]
) (
    // input logic[7:0][3:0] ports[8][10], my_grid,
    // a, b, c
);

input my_type_t[8:0][9:0] a[10][12];

output b;

logic[4:0] b[3];

endmodule